library verilog;
use verilog.vl_types.all;
entity IOTest_vlg_vec_tst is
end IOTest_vlg_vec_tst;
