module lcd_interface()

endmodule
