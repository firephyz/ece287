module MakeOutput(out);

	output [1:0] out;
	
	assign out = 2'b01;
	
endmodule
