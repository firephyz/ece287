library verilog;
use verilog.vl_types.all;
entity Lcd_vlg_vec_tst is
end Lcd_vlg_vec_tst;
