library verilog;
use verilog.vl_types.all;
entity lab_verilog_example_vlg_vec_tst is
end lab_verilog_example_vlg_vec_tst;
